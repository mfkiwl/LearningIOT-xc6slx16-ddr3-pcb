library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity uart is
    Port (tx:out BIT);
end uart;

architecture Behavioral of uart is

begin


end Behavioral;